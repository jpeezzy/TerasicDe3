
reg [512]abc[64]=
{
512'h6a09e667bb67ae853c6ef372a54ff53a510e527f9b05688c1f83d9ab5be0cd19,
512'h5d6aebcd6a09e667bb67ae853c6ef372fa2a4622510e527f9b05688c1f83d9ab,
512'h5a6ad9ad5d6aebcd6a09e667bb67ae8578ce7989fa2a4622510e527f9b05688c,
512'hc8c347a75a6ad9ad5d6aebcd6a09e667f92939eb78ce7989fa2a4622510e527f,
512'hd550f666c8c347a75a6ad9ad5d6aebcd24e00850f92939eb78ce7989fa2a4622,
512'h04409a6ad550f666c8c347a75a6ad9ad43ada24524e00850f92939eb78ce7989,
512'h2b4209f504409a6ad550f666c8c347a7714260ad43ada24524e00850f92939eb,
512'he50303802b4209f504409a6ad550f6669b27a401714260ad43ada24524e00850,
512'h85a07b5fe50303802b4209f504409a6a0c657a799b27a401714260ad43ada245,
512'h8e04ecb985a07b5fe50303802b4209f532ca2d8c0c657a799b27a401714260ad,
512'h8c87346b8e04ecb985a07b5fe50303801cc9259632ca2d8c0c657a799b27a401,
512'h4798a3f48c87346b8e04ecb985a07b5f436b23e81cc9259632ca2d8c0c657a79,
512'hf71fc5a94798a3f48c87346b8e04ecb9816fd6e9436b23e81cc9259632ca2d8c,
512'h87912990f71fc5a94798a3f48c87346b1e578218816fd6e9436b23e81cc92596,
512'hd932eb1687912990f71fc5a94798a3f4745a48de1e578218816fd6e9436b23e8,
512'hc0645fded932eb1687912990f71fc5a90b92f20c745a48de1e578218816fd6e9,
512'hb0fa238ec0645fded932eb168791299007590dcd0b92f20c745a48de1e578218,
512'h21da9a9bb0fa238ec0645fded932eb168034229c07590dcd0b92f20c745a48de,
512'hc2fbd9d121da9a9bb0fa238ec0645fde846ee4548034229c07590dcd0b92f20c,
512'hfe777bbfc2fbd9d121da9a9bb0fa238ecc899961846ee4548034229c07590dcd,
512'he1f20c33fe777bbfc2fbd9d121da9a9bb0638179cc899961846ee4548034229c,
512'h9dc68b63e1f20c33fe777bbfc2fbd9d18ada8930b0638179cc899961846ee454,
512'hc2606d6d9dc68b63e1f20c33fe777bbfe12579708ada8930b0638179cc899961,
512'ha7a3623fc2606d6d9dc68b63e1f20c3349f5114ae12579708ada8930b0638179,
512'hc5d53d8da7a3623fc2606d6d9dc68b63aa47c34749f5114ae12579708ada8930,
512'h1c2c2838c5d53d8da7a3623fc2606d6d2823ef91aa47c34749f5114ae1257970,
512'hcde8037d1c2c2838c5d53d8da7a3623f14383d8e2823ef91aa47c34749f5114a,
512'hb62ec4bccde8037d1c2c2838c5d53d8dc74c651614383d8e2823ef91aa47c347,
512'h77d37528b62ec4bccde8037d1c2c2838edffbff8c74c651614383d8e2823ef91,
512'h363482c977d37528b62ec4bccde8037d6112a3b7edffbff8c74c651614383d8e,
512'ha0060b30363482c977d37528b62ec4bcade794376112a3b7edffbff8c74c6516,
512'hea992a22a0060b30363482c977d375280109ab3aade794376112a3b7edffbff8,
512'h73b33bf5ea992a22a0060b30363482c9ba5911120109ab3aade794376112a3b7,
512'h98e1250773b33bf5ea992a22a0060b309cd9f5f6ba5911120109ab3aade79437,
512'hfe604df598e1250773b33bf5ea992a2259249dd39cd9f5f6ba5911120109ab3a,
512'ha9a7738cfe604df598e1250773b33bf5085f383359249dd39cd9f5f6ba591112,
512'h65a0cfe4a9a7738cfe604df598e12507f4b002d6085f383359249dd39cd9f5f6,
512'h41a65cb165a0cfe4a9a7738cfe604df50772a26bf4b002d6085f383359249dd3,
512'h34df160441a65cb165a0cfe4a9a7738ca507a53d0772a26bf4b002d6085f3833,
512'h6dc57a8a34df160441a65cb165a0cfe4f0781bc8a507a53d0772a26bf4b002d6,
512'h79ea687a6dc57a8a34df160441a65cb11efbc0a0f0781bc8a507a53d0772a26b,
512'hd667076679ea687a6dc57a8a34df160426352d631efbc0a0f0781bc8a507a53d,
512'hdf46652fd667076679ea687a6dc57a8a838b271126352d631efbc0a0f0781bc8,
512'h17aa0dfedf46652fd667076679ea687adecd4715838b271126352d631efbc0a0,
512'h9d4baf9317aa0dfedf46652fd6670766fda24c2edecd4715838b271126352d63,
512'h266288159d4baf9317aa0dfedf46652fa80f11f0fda24c2edecd4715838b2711,
512'h72ab4b91266288159d4baf9317aa0dfeb7755da1a80f11f0fda24c2edecd4715,
512'ha14c14b072ab4b91266288159d4baf93d57b94a9b7755da1a80f11f0fda24c2e,
512'h4172328da14c14b072ab4b9126628815fecf0bc6d57b94a9b7755da1a80f11f0,
512'h05757ceb4172328da14c14b072ab4b91bd714038fecf0bc6d57b94a9b7755da1,
512'hf11bfaa805757ceb4172328da14c14b06e5c390cbd714038fecf0bc6d57b94a9,
512'h7a0508a1f11bfaa805757ceb4172328d52f1ccf76e5c390cbd714038fecf0bc6,
512'h886e7a227a0508a1f11bfaa805757ceb49231c1e52f1ccf76e5c390cbd714038,
512'h101fd28f886e7a227a0508a1f11bfaa8529e7d0049231c1e52f1ccf76e5c390c,
512'hf5702fdb101fd28f886e7a227a0508a19f4787c3529e7d0049231c1e52f1ccf7,
512'h3ec45cdbf5702fdb101fd28f886e7a22e50e1b4f9f4787c3529e7d0049231c1e,
512'h38cc99133ec45cdbf5702fdb101fd28f54cb266be50e1b4f9f4787c3529e7d00,
512'hfcd1887b38cc99133ec45cdbf5702fdb9b5e906c54cb266be50e1b4f9f4787c3,
512'hc062d46ffcd1887b38cc99133ec45cdb7e44008e9b5e906c54cb266be50e1b4f,
512'hffb70472c062d46ffcd1887b38cc99136d83bfc67e44008e9b5e906c54cb266b,
512'hb6ae8fffffb70472c062d46ffcd1887bb21bad3d6d83bfc67e44008e9b5e906c,
512'hb85e2ce9b6ae8fffffb70472c062d46f961f4894b21bad3d6d83bfc67e44008e,
512'h04d24d6cb85e2ce9b6ae8fffffb70472948d25b6961f4894b21bad3d6d83bfc6,
512'hd39a216504d24d6cb85e2ce9b6ae8ffffb121210948d25b6961f4894b21bad3d,
512'h506e3058d39a216504d24d6cb85e2ce95ef50f24fb121210948d25b6961f4894
}
