`define sampleInput 512'h5105b8184c971573f8363c4d67abd3b87121d04a61c1a6cd16ff687c52aff4924159689767445b6046dd43d7c0aefdd2edd4bfd2fa1ef7e1ed93c97b1965a326

