//Here are all the constants 
`define h0 8'h6a09e667
`define h1 8'hbb67ae85
`define h2 8'h3c6ef372
`define h3 8'ha54ff53a
`define h4 8'h510e527f
`define h5 8'h9b05688c
`define h6 8'h1f83d9ab
`define h7 8'h5be0cd19

integer k[0:63] = {
8'h428a2f98, 8'h71374491, 8'hb5c0fbcf, 8'he9b5dba5, 8'h3956c25b, 
8'h59f111f1, 8'h923f82a4, 8'hab1c5ed5, 8'hd807aa98, 8'h12835b01, 
8'h243185be, 8'h550c7dc3, 8'h72be5d74, 8'h80deb1fe, 8'h9bdc06a7, 
8'hc19bf174, 8'he49b69c1, 8'hefbe4786, 8'h0fc19dc6, 8'h240ca1cc, 
8'h2de92c6f, 8'h4a7484aa, 8'h5cb0a9dc, 8'h76f988da, 8'h983e5152, 
8'ha831c66d, 8'hb00327c8, 8'hbf597fc7, 8'hc6e00bf3, 8'hd5a79147, 
8'h06ca6351, 8'h14292967, 8'h27b70a85, 8'h2e1b2138, 8'h4d2c6dfc, 
8'h53380d13, 8'h650a7354, 8'h766a0abb, 8'h81c2c92e, 8'h92722c85, 
8'ha2bfe8a1, 8'ha81a664b, 8'hc24b8b70, 8'hc76c51a3, 8'hd192e819, 
8'hd6990624, 8'hf40e3585, 8'h106aa070, 8'h19a4c116, 8'h1e376c08, 
8'h2748774c, 8'h34b0bcb5, 8'h391c0cb3, 8'h4ed8aa4a, 8'h5b9cca4f, 
8'h682e6ff3, 8'h748f82ee, 8'h78a5636f, 8'h84c87814, 8'h8cc70208, 
8'h90befffa, 8'ha4506ceb, 8'hbef9a3f7, 8'hc67178f2
};


